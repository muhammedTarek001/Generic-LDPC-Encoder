`ifndef BG2_pkg_PARAM
`define BG2_pkg_PARAM

package BG2_pkg;
  import LDPC_pkg::* ;




  parameter          BG2_MAX_TRANSFORMS      = 150;

  parameter bit[6:0] BG2_NON_MINUS_ONE_ELEMENTS [0:BG2_MAX_TRANSFORMS-1] = '{
0 ,1 ,2 ,3 ,6 ,9  ,

0 , 3 , 4 , 5 , 6 , 7 , 8 , 9  ,

0 , 1 , 3 , 4 , 8  ,

1 , 2 , 4 , 5 , 6 , 7 , 8 , 9  ,

0 , 1 , 11  ,

0 , 1 , 5 , 7 , 11  ,

0 , 5 , 7 , 9 , 11  ,

1 , 5 , 7 , 11 , 13  ,

0 , 1 , 12  ,

1 , 8 , 10 , 11  ,

0 , 1 , 6 , 7  ,

0 , 7 , 9 , 13  ,

1 , 3 , 11  ,

0 , 1 , 8 , 13  ,

1 , 6 , 11 , 13  ,

0 , 10 , 11  ,

1 , 9 , 11 , 12  ,

1 , 5 , 11 , 12  ,

0 , 6 , 7  ,

0 , 1 , 10  ,

1 , 4 , 11  ,

0 , 8 , 13  ,

1 , 2  ,

0 , 3 , 5  ,

1 , 2 , 9  ,

0 , 5  ,

2 , 7 , 12 , 13  ,

0 , 6  ,

1 , 2 , 5  ,

0 , 4  ,

2 , 5 , 7 , 9  ,

1 , 13  ,

0 , 5 , 12  ,

2 , 7 , 10  ,

0 , 12 , 13  ,

1 , 5 , 11  ,

0 , 2 , 7  ,

10 , 13  ,

1 , 5 , 11  ,

0 , 7 , 12  ,

2 , 10 , 13  ,

1 , 5 , 11
};







  parameter bit [8:0] BG2_ILS_0 [0:BG2_MAX_TRANSFORMS-1] = '{
9, 117, 204, 26, 189, 205, 
 
167, 166, 253, 125, 226, 156, 224, 252, 
 
81, 114, 44, 52, 240, 
 
8, 58, 158, 104, 209, 54, 18, 128, 
 
179, 214, 71, 
 
231, 41, 194, 159, 103, 
 
155, 228, 45, 28, 158, 
 
129, 147, 140, 3, 116, 
 
142, 94, 230, 
 
203, 205, 61, 247, 
 
11, 185, 0, 117, 
 
11, 236, 210, 56, 
 
63, 111, 14, 
 
83, 2, 38, 222, 
 
115, 145, 3, 232, 
 
51, 175, 213, 
 
203, 142, 8, 242, 
 
254, 124, 114, 64, 
 
220, 194, 50, 
 
87, 20, 185, 
 
26, 105, 29, 
 
76, 42, 210, 
 
222, 63, 
 
23, 235, 238, 
 
46, 139, 8, 
 
228, 156, 
 
29, 143, 160, 122, 
 
8, 151, 
 
98, 101, 135, 
 
18, 28, 
 
71, 240, 9, 84, 
 
106, 1, 
 
242, 44, 166, 
 
132, 164, 235, 
 
147, 85, 36, 
 
57, 40, 63, 
 
140, 38, 154, 
 
219, 151, 
 
31, 66, 38, 
 
239, 172, 34, 
 
0, 75, 120, 
 
129, 229, 118
  };








  parameter bit [8:0] BG2_ILS_1 [0:BG2_MAX_TRANSFORMS-1] = '{
174, 97, 166, 66, 71, 172, 
 
27, 36, 48, 92, 31, 187, 185, 3, 
 
25, 114, 117, 110, 114, 
 
136, 175, 113, 72, 123, 118, 28, 186, 
 
72, 74, 29, 
 
10, 44, 121, 80, 48, 
 
129, 92, 100, 49, 184, 
 
80, 186, 16, 102, 143, 
 
118, 70, 152, 
 
28, 132, 185, 178, 
 
59, 104, 22, 52, 
 
32, 92, 174, 154, 
 
39, 93, 11, 
 
49, 125, 35, 166, 
 
19, 118, 21, 163, 
 
68, 63, 81, 
 
87, 177, 135, 64, 
 
158, 23, 9, 6, 
 
186, 6, 46, 
 
58, 42, 156, 
 
76, 61, 153, 
 
157, 175, 67, 
 
20, 52, 
 
106, 86, 95, 
 
182, 153, 64, 
 
45, 21, 
 
67, 137, 55, 85, 
 
103, 50, 
 
70, 111, 168, 
 
110, 17, 
 
120, 154, 52, 56, 
 
3, 170, 
 
84, 8, 17, 
 
165, 179, 124, 
 
173, 177, 12, 
 
77, 184, 18, 
 
25, 151, 170, 
 
37, 31, 
 
84, 151, 190, 
 
93, 132, 57, 
 
103, 107, 163, 
 
147, 7, 60
  };
  






  parameter bit [8:0] BG2_ILS_2 [0:BG2_MAX_TRANSFORMS-1] = '{
0, 0, 0, 0, 0, 0, 
 
137, 124, 0, 0, 88, 0, 0, 55, 
 
20, 94, 99, 9, 108, 
 
38, 15, 102, 146, 12, 57, 53, 46, 
 
0, 136, 157, 
 
0, 131, 142, 141, 64, 
 
0, 124, 99, 45, 148, 
 
0, 45, 148, 96, 78, 
 
0, 65, 87, 
 
0, 97, 51, 85, 
 
0, 17, 156, 20, 
 
0, 7, 4, 2, 
 
0, 113, 48, 
 
0, 112, 102, 26, 
 
0, 138, 57, 27, 
 
0, 73, 99, 
 
0, 79, 111, 143, 
 
0, 24, 109, 18, 
 
0, 18, 86, 
 
0, 158, 154, 
 
0, 148, 104, 
 
0, 17, 33, 
 
0, 4, 
 
0, 75, 158, 
 
0, 69, 87, 
 
0, 65, 
 
0, 100, 13, 7, 
 
0, 32, 
 
0, 126, 110, 
 
0, 154, 
 
0, 35, 51, 134, 
 
0, 20, 
 
0, 20, 122, 
 
0, 88, 13, 
 
0, 19, 78, 
 
0, 157, 6, 
 
0, 63, 82, 
 
0, 144, 
 
0, 93, 19, 
 
0, 24, 138, 
 
0, 36, 143, 
 
0, 2, 55
  };
  






  parameter bit [8:0] BG2_ILS_3 [0:BG2_MAX_TRANSFORMS-1] = '{
72, 110, 23, 181, 95, 8, 
 
53, 156, 115, 156, 115, 200, 29, 31, 
 
152, 131, 46, 191, 91, 
 
185, 6, 36, 124, 124, 110, 156, 133, 
 
200, 16, 101, 
 
185, 138, 170, 219, 193, 
 
123, 55, 31, 222, 209, 
 
103, 13, 105, 150, 181, 
 
147, 43, 152, 
 
2, 30, 184, 83, 
 
174, 150, 8, 56, 
 
99, 138, 110, 99, 
 
46, 217, 109, 
 
37, 113, 143, 140, 
 
36, 95, 40, 116, 
 
116, 200, 110, 
 
75, 158, 134, 97, 
 
48, 132, 206, 2, 
 
68, 16, 156, 
 
35, 138, 86, 
 
6, 20, 141, 
 
80, 43, 81, 
 
49, 1, 
 
156, 54, 134, 
 
153, 88, 63, 
 
211, 94, 
 
90, 6, 221, 6, 
 
27, 118, 
 
216, 212, 193, 
 
108, 61, 
 
106, 44, 185, 176, 
 
147, 182, 
 
108, 21, 110, 
 
71, 12, 109, 
 
29, 201, 69, 
 
91, 165, 55, 
 
1, 175, 83, 
 
40, 12, 
 
37, 97, 46, 
 
106, 181, 154, 
 
98, 35, 36, 
 
120, 101, 81
  };






  parameter bit [8:0] BG2_ILS_4 [0:BG2_MAX_TRANSFORMS-1] = '{
3, 26, 53, 35, 115, 127, 
 
19, 94, 104, 66, 84, 98, 69, 50, 
 
95, 106, 92, 110, 111, 
 
120, 121, 22, 4, 73, 49, 128, 79, 
 
42, 24, 51, 
 
40, 140, 84, 137, 71, 
 
109, 87, 107, 133, 139, 
 
97, 135, 35, 108, 65, 
 
70, 69, 88, 
 
97, 40, 24, 49, 
 
46, 41, 101, 96, 
 
28, 30, 116, 64, 
 
33, 122, 131, 
 
76, 37, 62, 47, 
 
143, 51, 130, 97, 
 
139, 96, 128, 
 
48, 9, 28, 8, 
 
120, 43, 65, 42, 
 
17, 106, 142, 
 
79, 28, 41, 
 
2, 103, 78, 
 
91, 75, 81, 
 
54, 132, 
 
68, 115, 56, 
 
30, 42, 101, 
 
128, 63, 
 
142, 28, 100, 133, 
 
13, 10, 
 
106, 77, 43, 
 
133, 25, 
 
87, 56, 104, 70, 
 
80, 139, 
 
32, 89, 71, 
 
135, 6, 2, 
 
37, 25, 114, 
 
60, 137, 93, 
 
121, 129, 26, 
 
97, 56, 
 
1, 70, 1, 
 
119, 32, 142, 
 
6, 73, 102, 
 
48, 47, 19
  };
  






  parameter bit [8:0] BG2_ILS_5 [0:BG2_MAX_TRANSFORMS-1] = '{
156, 143, 14, 3, 40, 123, 
 
17, 65, 63, 1, 55, 37, 171, 133, 
 
98, 168, 107, 82, 142, 
 
53, 174, 174, 127, 17, 89, 17, 105, 
 
86, 67, 83, 
 
79, 84, 35, 103, 60, 
 
47, 154, 10, 155, 29, 
 
48, 125, 24, 47, 55, 
 
53, 31, 161, 
 
104, 142, 99, 64, 
 
111, 25, 174, 23, 
 
91, 175, 24, 141, 
 
122, 11, 4, 
 
29, 91, 27, 127, 
 
11, 145, 8, 166, 
 
137, 103, 40, 
 
78, 158, 17, 165, 
 
134, 23, 62, 163, 
 
173, 31, 22, 
 
13, 135, 145, 
 
128, 52, 173, 
 
156, 166, 40, 
 
18, 163, 
 
110, 132, 150, 
 
113, 108, 61, 
 
72, 136, 
 
36, 38, 53, 145, 
 
42, 104, 
 
64, 24, 149, 
 
139, 161, 
 
84, 173, 93, 29, 
 
117, 148, 
 
116, 73, 142, 
 
105, 137, 29, 
 
11, 41, 162, 
 
126, 152, 172, 
 
73, 154, 129, 
 
167, 38, 
 
112, 7, 19, 
 
109, 6, 105, 
 
160, 156, 82, 
 
132, 6, 8
  };
  






  parameter bit [8:0] BG2_ILS_6 [0:BG2_MAX_TRANSFORMS-1] = '{
143, 19, 176, 165, 196, 13, 
 
18, 27, 3, 102, 185, 17, 14, 180, 
 
126, 163, 47, 183, 132, 
 
36, 48, 18, 111, 203, 3, 191, 160, 
 
43, 27, 117, 
 
136, 49, 36, 132, 62, 
 
7, 34, 198, 168, 12, 
 
163, 78, 143, 107, 58, 
 
101, 177, 22, 
 
186, 27, 205, 81, 
 
125, 60, 177, 51, 
 
39, 29, 35, 8, 
 
18, 155, 49, 
 
32, 53, 95, 186, 
 
91, 20, 52, 109, 
 
174, 108, 102, 
 
125, 31, 54, 176, 
 
57, 201, 142, 35, 
 
129, 203, 140, 
 
110, 124, 52, 
 
196, 35, 114, 
 
10, 122, 23, 
 
202, 126, 
 
52, 170, 13, 
 
113, 161, 88, 
 
197, 194, 
 
164, 172, 49, 161, 
 
168, 193, 
 
14, 186, 46, 
 
50, 27, 
 
70, 17, 50, 6, 
 
115, 189, 
 
110, 0, 163, 
 
163, 173, 179, 
 
197, 191, 193, 
 
157, 167, 181, 
 
197, 167, 179, 
 
181, 193, 
 
157, 173, 191, 
 
181, 157, 173, 
 
193, 163, 179, 
 
191, 197, 167
  };






  parameter bit [8:0] BG2_ILS_7 [0:BG2_MAX_TRANSFORMS-1] = '{
145, 131, 71, 21, 23, 112, 
 
142, 174, 183, 27, 96, 23, 9, 167, 
 
74, 31, 3, 53, 155, 
 
239, 171, 95, 110, 159, 199, 43, 75, 
 
29, 140, 180, 
 
121, 41, 169, 88, 207, 
 
137, 72, 172, 124, 56, 
 
86, 186, 87, 172, 154, 
 
176, 169, 225, 
 
167, 238, 48, 68, 
 
38, 217, 208, 232, 
 
178, 214, 168, 51, 
 
124, 122, 72, 
 
48, 57, 167, 219, 
 
82, 232, 204, 162, 
 
38, 217, 157, 
 
170, 23, 175, 202, 
 
196, 173, 195, 218, 
 
128, 211, 210, 
 
39, 84, 88, 
 
117, 227, 6, 
 
238, 13, 11, 
 
195, 44, 
 
5, 94, 111, 
 
81, 19, 130, 
 
66, 95, 
 
146, 66, 190, 86, 
 
64, 181, 
 
7, 144, 16, 
 
25, 57, 
 
37, 139, 221, 17, 
 
201, 46, 
 
179, 14, 116, 
 
46, 2, 106, 
 
184, 135, 141, 
 
85, 225, 175, 
 
178, 112, 106, 
 
154, 114, 
 
42, 41, 105, 
 
167, 45, 189, 
 
78, 67, 180, 
 
53, 215, 230
  };



endpackage

`endif