`ifndef BG1_pkg_PARAM
`define BG1_pkg_PARAM

package BG1_pkg;
  import LDPC_pkg::* ;
  

parameter     BG1_MAX_TRANSFORMS      = 265;

parameter bit[5:0] BG1_NON_MINUS_ONE_ELEMENTS [0:BG1_MAX_TRANSFORMS-1] = '{
0 ,1 ,2 ,3 ,5 ,6 ,9 ,10,11,12,13,15,16,18,19,20,21,

0 ,2 ,3 ,4 ,5 ,7 ,8 ,9 ,11,12,14,15,16,17,19,21,

0 ,1 ,2 ,4 ,5 ,6 ,7 ,8 ,9 ,10,13,14,15,17,18,19,20,

0 ,1 ,3 ,4 ,6 ,7 ,8 ,10,11,12,13,14,16,17,18,20,21,

0,1,

0,1,3,12,16,21,22,

0 ,6 ,10,11,13,17,18,20,

0 ,1 ,4 ,7 ,8 ,14,

0 ,1 ,3 ,12 ,16 ,19 ,21 ,22 ,24 ,

0 ,1 ,10 ,11 ,13 ,17 ,18 ,20 ,

1 ,2 ,4 ,7 ,8 ,14 ,

0 ,1 ,12 ,16 ,21 ,22 ,23 ,

0 , 1 , 10 , 11 , 13 , 18 ,

0 , 3 , 7 , 20 , 23 ,

0 , 12 , 15 , 16 , 17 , 21 ,

0 , 1 , 10 , 13 , 18 , 25 ,

1 , 3 , 11 , 20 , 22 ,

0 , 14 , 16 , 17 , 21 ,

1 , 12 , 13 , 18 , 19 ,

0 , 1 , 7 , 8 , 10 ,

0 , 3 , 9 , 11 , 22 ,

1 , 5 , 16 , 20 , 21 ,

0 , 12 , 13 , 17 ,

1 , 2 , 10 , 18 ,

0 , 3 , 4 , 11 , 22 ,

1 , 6 , 7 , 14 ,

0 , 2 , 4 , 15 ,

1 , 6 , 8 ,

0 , 4 , 19 , 21 ,

1 , 14 , 18 , 25 ,

0 , 10 , 13 , 24 ,

1 , 7 , 22 , 25 ,

0 , 12 , 14 , 24 ,

1 , 2 , 11 , 21 ,

0 , 7 , 15 , 17 ,

1 , 6 , 12 , 22 ,

0 , 14 , 15 , 18 ,

1 , 13 , 23 ,

0 , 9 , 10 , 12 ,

1 , 3 , 7 , 19 ,

0 , 8 , 17 ,

1 , 3 , 9 , 18 ,

0 , 4 , 24 ,

1 , 16 , 18 , 25 ,

0 , 7 , 9 , 22 ,

1 , 6 , 10
};



  parameter bit [8:0] BG1_ILS_0 [0:BG1_MAX_TRANSFORMS-1] = '{
250,69,226,159,100,10,59,229,110,191,9,195,23,190,35,239,31,
 
2,239,117,124,71,222,104,173,220,102,109,132,142,155,255,28,
 
106,111,185,63,117,93,229,177,95,39,142,225,225,245,205,251,117,
 
121,89,84,20,150,131,243,136,86,246,219,211,240,76,244,144,12,
 
157,102,
 
205,236,194,231,28,123,115,
 
183,22,28,67,244,11,157,211,
 
220,44,159,31,167,104,
 
112,4,7,211,102,164,109,241,90,
 
103,182,109,21,142,14,61,216,
 
98,149,167,160,49,58,
 
77,41,83,182,78,252,22,
 
160,42,21,32,234,7,
 
177,248,151,185,62,
 
206,55,206,127,16,229,
 
40,96,65,63,75,179,
 
64,49,49,51,154,
 
7,164,59,1,144,
 
42,233,8,155,147,
 
60,73,72,127,224,
 
151,186,217,47,160,
 
249,121,109,131,171,
 
64,142,188,158,
 
156,147,170,152,
 
112,86,236,116,222,
 
23,136,116,182,
 
195,243,215,61,
 
25,104,194,
 
128,165,181,63,
 
86,236,84,6,
 
216,73,120,9,
 
95,177,172,61,
 
221,112,199,121,
 
2,187,41,211,
 
127,167,164,159,
 
161,197,207,103,
 
37,105,51,120,
 
198,220,122,
 
167,151,157,163,
 
173,139,149,0,
 
157,137,149,
 
167,173,139,151,
 
149,157,137,
 
151,163,173,139,
 
139,157,163,173,
 
149,151,167
}; 





























  parameter bit [8:0] BG1_ILS_1 [0:BG1_MAX_TRANSFORMS-1] = '{
307,19,50,369,181,216,317,288,109,17,357,215,106,242,180,330,346,
 
76,76,73,288,144,331,331,178,295,342,217,99,354,114,331,112,
 
205,250,328,332,256,161,267,160,63,129,200,88,53,131,240,205,13,
 
276,87,0,275,199,153,56,132,305,231,341,212,304,300,271,39,357,
 
332,181,
 
195,14,115,166,241,51,157,
 
278,257,1,351,92,253,18,225,
 
9,62,316,333,290,114,
 
307,179,165,18,39,224,368,67,170,
 
366,232,321,133,57,303,63,82,
 
101,339,274,111,383,354,
 
48,102,8,47,188,334,115,
 
77,186,174,232,50,74,
 
313,177,266,115,370,
 
142,248,137,89,347,12,
 
241,2,210,318,55,269,
 
13,338,57,289,57,
 
260,303,81,358,375,
 
130,163,280,132,4,
 
145,213,344,242,197,
 
187,206,264,341,59,
 
205,102,328,213,97,
 
30,11,233,22,
 
24,89,61,27,
 
298,158,235,339,234,
 
72,17,383,312,
 
71,81,76,136,
 
194,194,101,
 
222,19,244,274,
 
252,5,147,78,
 
159,229,260,90,
 
100,215,258,256,
 
102,201,175,287,
 
323,8,361,105,
 
230,148,202,312,
 
320,335,2,266,
 
210,313,297,21,
 
269,82,115,
 
185,177,289,214,
 
258,93,346,297,
 
175,37,312,
 
52,314,139,288,
 
113,14,218,
 
113,132,114,168,
 
80,78,163,274,
 
135,149,15
  };

















  parameter bit [8:0] BG1_ILS_2 [0:BG1_MAX_TRANSFORMS-1] = '{
73,15,103,49,240,39,15,162,215,164,133,298,110,113,16,189,32,
 
303,294,27,261,161,133,4,80,129,300,76,266,72,83,260,301,
 
68,7,80,280,38,227,202,200,71,106,295,283,301,184,246,230,276,
 
220,208,30,197,61,175,79,281,303,253,164,53,44,28,77,319,68,
 
233,205,
 
83,292,50,318,201,267,279,
 
289,21,293,13,232,302,138,235,
 
12,88,207,50,25,76,
 
295,133,130,231,296,110,269,245,154,
 
189,244,36,286,151,267,135,209,
 
14,80,211,75,161,311,
 
16,147,290,289,177,43,280,
 
229,235,169,48,105,52,
 
39,302,303,160,37,
 
78,299,54,61,179,258,
 
229,290,60,130,184,51,
 
69,140,45,115,300,
 
257,147,128,51,228,
 
260,294,291,141,295,
 
64,181,101,270,41,
 
301,162,40,130,10,
 
79,175,132,283,103,
 
177,20,55,316,
 
249,50,133,105,
 
289,280,110,187,281,
 
172,295,96,46,
 
270,110,318,67,
 
210,29,304,
 
11,293,50,234,
 
27,308,117,29,
 
91,23,105,135,
 
222,308,66,162,
 
210,22,271,217,
 
170,20,140,33,
 
187,296,5,44,
 
207,158,55,285,
 
259,179,178,160,
 
298,15,115,
 
151,179,64,181,
 
102,77,192,208,
 
32,80,197,
 
154,47,124,207,
 
226,65,126,
 
228,69,176,102,
 
234,227,259,260,
 
101,228,126
  };










    parameter bit [8:0] BG1_ILS_3 [0:BG1_MAX_TRANSFORMS-1] = '{
223,16,94,91,74,10,0,205,216,21,215,14,70,141,198,104,81,
 
141,45,151,46,119,157,133,87,206,93,79,9,118,194,31,187,
 
207,203,31,176,180,186,95,153,177,70,77,214,77,198,117,223,90,
 
201,18,165,5,45,142,16,34,155,213,147,69,96,74,99,30,158,
 
170,10,
 
164,59,86,80,182,130,153,
 
158,119,113,21,63,51,136,116,
 
17,76,104,100,150,158,
 
33,95,4,217,204,39,58,44,201,
 
9,37,213,105,89,185,109,218,
 
82,165,174,19,194,103,
 
52,11,2,35,32,84,201,
 
142,175,136,3,28,182,
 
81,56,72,217,78,
 
14,175,211,191,51,43,
 
90,120,131,209,209,81,
 
154,164,43,189,101,
 
56,110,200,63,4,
 
199,110,200,143,186,
 
8,6,103,198,8,
 
105,210,121,214,183,
 
192,131,220,50,106,
 
53,0,3,148,
 
88,203,168,122,
 
49,157,64,193,124,
 
1,166,65,81,
 
107,176,212,127,
 
208,141,174,
 
146,153,217,114,
 
150,11,53,68,
 
34,130,210,123,
 
175,49,177,128,
 
192,209,58,30,
 
114,49,161,137,
 
82,186,68,150,
 
192,173,26,187,
 
222,157,0,6,
 
81,195,138,
 
123,90,73,10,
 
12,77,49,114,
 
67,45,96,
 
23,215,60,167,
 
114,91,78,
 
206,22,134,161,
 
84,4,9,12,
 
184,121,29
  };





  parameter bit [8:0] BG1_ILS_4 [0:BG1_MAX_TRANSFORMS-1] = '{
211,198,188,186,219,4,29,144,116,216,115,233,144,95,216,73,261,
 
179,162,223,256,160,76,202,117,109,15,72,152,158,147,156,119,
 
258,167,220,133,243,202,218,63,0,3,74,229,0,216,269,200,234,
 
187,145,166,108,82,132,197,41,162,57,36,115,242,165,0,113,108,
 
246,235,
 
261,181,72,283,254,79,144,
 
80,144,169,90,59,177,151,108,
 
169,189,154,184,104,164,
 
54,0,252,41,98,46,15,230,54,
 
162,159,93,134,45,132,76,209,
 
178,1,28,267,234,201,
 
55,23,274,181,273,39,26,
 
225,162,244,151,238,243,
 
231,0,216,47,36,
 
0,186,253,16,0,79,
 
170,0,183,108,68,64,
 
270,13,99,54,0,
 
153,137,0,0,162,
 
161,151,0,241,144,
 
0,0,118,144,0,
 
265,81,90,144,228,
 
64,46,266,9,18,
 
72,189,72,257,
 
180,0,0,165,
 
236,199,0,266,0,
 
205,0,0,183,
 
0,0,0,277,
 
45,36,72,
 
275,0,155,62,
 
0,180,0,42,
 
0,90,252,173,
 
144,144,166,19,
 
0,211,36,162,
 
0,0,76,18,
 
197,0,108,0,
 
199,278,0,205,
 
216,16,0,0,
 
72,144,0,
 
190,0,0,0,
 
153,0,165,117,
 
216,144,2,
 
0,0,0,183,
 
27,0,35,
 
52,243,0,270,
 
18,0,0,57,
 
168,0,144
};











  parameter bit [8:0] BG1_ILS_5 [0:BG1_MAX_TRANSFORMS-1] = '{
294,118,167,330,207,165,243,250,1,339,201,53,347,304,167,47,188,
 
77,225,96,338,268,112,302,50,167,253,334,242,257,133,9,302,
 
226,35,213,302,111,265,128,237,294,127,110,286,125,131,163,210,7,
 
97,94,49,279,139,166,91,106,246,345,269,185,249,215,143,121,121,
 
42,256,
 
219,130,251,322,295,258,283,
 
294,73,330,99,172,150,284,305,
 
3,103,224,297,215,39,
 
348,75,22,312,224,17,59,314,244,
 
156,88,293,111,92,152,23,337,
 
175,253,27,231,49,267,
 
25,322,200,351,166,338,192,
 
123,217,142,110,176,76,
 
311,251,265,94,81,
 
22,322,277,156,66,78,
 
176,348,15,81,176,113,
 
190,293,332,331,114,
 
110,228,247,116,190,
 
47,286,246,181,73,
 
87,110,147,258,204,
 
89,65,155,244,30,
 
162,264,346,143,109,
 
280,157,236,113,
 
18,6,181,304,
 
38,170,249,288,194,
 
279,255,111,54,
 
325,326,226,99,
 
91,326,268,
 
102,1,40,167,
 
273,104,243,107,
 
171,16,95,212,
 
101,297,279,222,
 
351,265,338,83,
 
56,304,141,101,
 
60,320,112,54,
 
100,210,195,268,
 
135,15,35,188,
 
319,236,85,
 
164,196,209,246,
 
236,264,37,272,
 
304,237,135,
 
123,77,25,272,
 
288,83,17,
 
210,3,53,167,
 
79,244,293,272,
 
82,67,235
};











  parameter bit [8:0] BG1_ILS_6 [0:BG1_MAX_TRANSFORMS-1] = '{
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
 
22,11,124,0,10,0,0,2,16,60,0,6,30,0,168,31,
 
132,37,21,180,4,149,48,38,122,195,155,28,85,47,179,42,66,
 
4,6,33,113,49,21,6,151,83,154,87,5,92,173,120,2,142,
 
24,204,
 
185,100,24,65,207,161,72,
 
6,27,163,50,48,24,38,91,
 
145,88,112,153,159,76,
 
172,2,131,141,96,99,101,35,116,
 
6,10,145,53,201,4,164,173,
 
126,77,156,16,12,70,
 
184,194,123,16,104,109,124,
 
6,20,203,153,104,207,
 
52,147,1,16,46,
 
1,202,118,130,1,2,
 
173,6,81,182,53,46,
 
88,198,160,122,182,
 
91,184,30,3,155,
 
1,41,167,68,148,
 
12,6,166,184,191,
 
6,12,15,5,30,
 
6,86,96,42,199,
 
44,58,130,131,
 
45,18,132,100,
 
9,125,191,28,6,
 
4,74,16,28,
 
21,142,192,197,
 
98,140,22,
 
4,1,40,93,
 
92,136,106,6,
 
2,88,112,20,
 
4,49,125,194,
 
6,126,63,20,
 
10,30,6,92,
 
4,153,197,155,
 
4,45,168,185,
 
6,200,177,43,
 
82,2,135,
 
91,64,198,100,
 
4,28,109,188,
 
10,84,12,
 
2,75,142,128,
 
163,10,162,
 
1,163,99,98,
 
4,6,142,3,
 
181,45,153
};








  parameter bit [8:0] BG1_ILS_7 [0:BG1_MAX_TRANSFORMS-1] = '{
135,227,126,134,84,83,53,225,205,128,75,135,217,220,90,105,137,
 
96,236,136,221,128,92,172,56,11,189,95,85,153,87,163,216,
 
189,4,225,151,236,117,179,92,24,68,6,101,33,96,125,67,230,
 
128,23,162,220,43,186,96,1,216,22,24,167,200,32,235,172,219,
 
64,211,
 
2,171,47,143,210,180,180,
 
199,22,23,100,92,207,52,13,
 
77,146,209,32,166,18,
 
181,105,141,223,177,145,199,153,38,
 
169,12,206,221,17,212,92,205,
 
116,151,70,230,115,84,
 
45,115,134,1,152,165,107,
 
186,215,124,180,98,80,
 
220,185,154,178,150,
 
124,144,182,95,72,76,
 
39,138,220,173,142,49,
 
78,152,84,5,205,
 
183,112,106,219,129,
 
183,215,180,143,14,
 
179,108,159,138,196,
 
77,187,203,167,130,
 
197,122,215,65,216,
 
25,47,126,178,
 
185,127,117,199,
 
32,178,2,156,58,
 
27,141,11,181,
 
163,131,169,98,
 
165,232,9,
 
32,43,200,205,
 
232,32,118,103,
 
170,199,26,105,
 
73,149,175,108,
 
103,110,151,211,
 
199,132,172,65,
 
161,237,142,180,
 
231,174,145,100,
 
11,207,42,100,
 
59,204,161,
 
121,90,26,140,
 
115,188,168,52,
 
4,103,30,
 
53,189,215,24,
 
222,170,71,
 
22,127,49,125,
 
191,211,187,148,
 
177,114,93
};



//::--------------------------------------------------------------------------------------------------------------------------------:://
//::--------------------------------------------------------------------------------------------------------------------------------:://



endpackage

`endif